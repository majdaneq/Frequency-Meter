-------------------------------------------------------------------------------
--
-- Title       : Fub3
-- Design      : Miernik_czestotliwosci
-- Author      : szymonbortel8@gmail.com
-- Company     : agh
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\szymo\Desktop\PSC_Projekt\miernik_czest\Miernik_czestotliwosci\src\Fub3.vhd
-- Generated   : Tue Jan 16 21:39:25 2018
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Fub3} architecture {Fub3}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Fub3 is
end Fub3;

--}} End of automatically maintained section

architecture Fub3 of Fub3 is
begin

	 -- enter your statements here --

end Fub3;
